library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

--This module acts as a buffer to save the data created by the renderer before
--it is written to the RAM. It holds data for eight pixel. The data is stored 
--in three shift registers (one for each colour). The bits are right shifted in 
--the registers. So the first rendered bit will be the LSB when the buffer is 
--full. A counter controls if the buffer is full. If so an output signal is set 
--to signalise that the buffer content needs to be written to the RAM. The 
--shift operation of the buffer can be activated with an external signal.
--There is no need to reset the buffer after writing its content to the RAM 
--because the internal counter is set to 0 when the next new data arrives and 
--the old content of the shift registers is replaced with the new data.

entity render_buffer is
  --ports:
  --clk             : system clock
  --reset           : synchronous reset
  --
  --i_shift_enable  : enable signal for the shift operation
  --i_rgb           : data vector for one pixel MSB(RRRGGGBB)LSB
  --
  --o_buffer_full   : signalises that the buffer is full
  --o_rgb_data : output for 32 pixel
  port (clk   : in std_logic := '0';
        reset : in std_logic := '0';

        i_shift_enable : in std_logic                     := '0';
        i_rgb          : in std_logic_vector (7 downto 0) := (others => '0');

        o_buffer_full : out std_logic                          := '1';
        o_rgb_data   : out std_logic_vector(32*8-1 downto 0) := (others => '0'));
--         o_red_data : out std_logic_vector (9 downto 0) := (others => '0');
--         o_green_data : out std_logic_vector (9 downto 0) := (others => '0');
--         o_blue_data : out std_logic_vector (9 downto 0) := (others => '0'));
end render_buffer;



architecture rtl of render_buffer is

--The following three signals store the content of the shift registers for the 
--three colours
  signal sr_rgb_data   : std_logic_vector (32*8-1 downto 0) := (others => '0');
--Counter for the number of bits already shifted to the registers.
  signal cnt_data      : integer range 0 to 31          := 0;

begin
  --Type : registered
  --Description : This buffer stores the data generated by the renderer. When 
  --    enabled the new data is shifted in the registers and the data counter 
  --    is increased to indicate how much data has already been stored in the 
  --    buffer and when it is full.
  process (clk)
  begin
    if (clk'event and clk = '1') then
      --Synchronous reset
      if (reset = '1') then
        sr_rgb_data   <= (others => '0');
        cnt_data      <= 0;
      --If shifting is enabled the new data is fed to the MSB of the shift 
      --register after a right shift was performed.
      elsif (i_shift_enable = '1') then
        sr_rgb_data   <= i_rgb & sr_rgb_data(32*8-1 downto 8);
        --If the counter has reached its maximum it is reset to 0.
        if (cnt_data = 31) then
          cnt_data <= 0;
        --The counter is increased by 1.
        else
          cnt_data <= cnt_data + 1;
        end if;
      end if;
    end if;
  end process;

  --The buffer full output is set when the data counter reaches 7 (one cycle 
  --before the buffer is full because it takes one clock cycle for the rnderer 
  --to react and stop rendering new data).
  o_buffer_full <= '1' when (cnt_data = 31)
                   else '0';
  --The content of the shift registers is assigned to the corresponding 
  --outputs.
  o_rgb_data   <= sr_rgb_data;
  
end rtl;

