library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity comb_logic is
   port (i_a : in std_logic := '0';
         i_b : in std_logic := '0';
         
         o_c : out std_logic := '0');
end comb_logic;


architecture rtl of comb_logic is
--signal declaration

  
begin





  
end rtl;
