library IEEE;
use IEEE.STD_LOGIC_1164.all;
use IEEE.NUMERIC_STD.all;

entity seq_logic is
  port (clk   : in std_logic := '0';
        reset : in std_logic := '0';

        i_a : in std_logic := '0';
        i_b : in std_logic := '0';

        o_q : out std_logic := '0');
end seq_logic;



architecture rtl of seq_logic is

-- signal declaration


-- component declaration


 
  
begin

-- component instantiation
 




end rtl;

