library verilog;
use verilog.vl_types.all;
entity cellram is
    generic(
        tACLK           : real    := 7.000000;
        tAPA            : real    := 20.000000;
        tAW             : real    := 70.000000;
        tBW             : real    := 70.000000;
        tCBPH           : real    := 5.000000;
        tCLK            : real    := 9.620000;
        tCSP            : real    := 3.000000;
        tCW             : real    := 70.000000;
        tHD             : real    := 2.000000;
        tKP             : real    := 3.000000;
        tPC             : real    := 20.000000;
        tRC             : real    := 70.000000;
        tSP             : real    := 3.000000;
        tVP             : real    := 5.000000;
        tVS             : real    := 70.000000;
        tWC             : real    := 70.000000;
        tWP             : real    := 45.000000;
        tAS             : real    := 0.000000;
        tAVH            : real    := 2.000000;
        tAVS            : real    := 5.000000;
        tCPH            : real    := 5.000000;
        tCVS            : real    := 7.000000;
        tDH             : real    := 0.000000;
        tDPDX           : real    := 10000.000000;
        tDW             : real    := 20.000000;
        tOW             : real    := 5.000000;
        tPU             : real    := 150000.000000;
        tVPH            : real    := 0.000000;
        tWPH            : real    := 10.000000;
        tWR             : real    := 0.000000;
        ADQ_BITS        : integer := 23;
        DQ_BITS         : integer := 16;
        BY_BITS         : integer := 2;
        ADDR_BITS       : integer := 23;
        COL_BITS        : integer := 7;
        MEM_BITS        : integer := 10;
        BCR             : integer := 2;
        RCR             : integer := 0;
        DIDR            : integer := 1;
        REG_SEL         : integer := 18;
        CR10            : integer := 1;
        CR15            : integer := 2;
        CR20            : integer := 3;
        GENERATION      : integer := 2;
        CR20WAIT_POLARITY: integer := 1;
        CRE_READ        : integer := 1;
        BCR_MASK        : integer := 261439;
        BCR_DEFAULT     : integer := 40223;
        RCR_MASK        : integer := 196759;
        RCR_DEFAULT     : integer := 16;
        DIDR_MASK       : integer := 262143;
        DIDR_DEFAULT    : integer := 835;
        DEBUG           : integer := 1;
        IDLE            : integer := 0;
        WR              : integer := 1;
        RD              : integer := 2;
        CFG_RD          : integer := 3;
        CFG_WR          : integer := 4
    );
    port(
        clk             : in     vl_logic;
        adv_n           : in     vl_logic;
        cre             : in     vl_logic;
        o_wait          : out    vl_logic;
        ce_n            : in     vl_logic;
        oe_n            : in     vl_logic;
        we_n            : in     vl_logic;
        lb_n            : in     vl_logic;
        ub_n            : in     vl_logic;
        addr            : in     vl_logic_vector;
        dq              : inout  vl_logic_vector
    );
end cellram;
